//
//
//

`define MINIMIG_ALTERA
//`define MINIMIG_XILINX
